// Erro semântico na linha 4: variável var1 já possui um valor.

var1 = var2 & var3
var1 = var2 | var3