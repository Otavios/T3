// Linha 3: @ - simbolo nao identificado

S = A ^ @B // xor
C = A & B // and